// AND Gate - Gate Level Modeling

module and_gate_gate_level(
    input a,
    input b,
    output y
);

and (y, a, b);

endmodule
